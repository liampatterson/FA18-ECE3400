`define SCREEN_WIDTH 176
`define SCREEN_HEIGHT 144
`define NUM_BARS 3
`define BAR_HEIGHT 48

module IMAGE_PROCESSOR (
	PIXEL_IN,
	CLK,
	VGA_PIXEL_X,
	VGA_PIXEL_Y,
	VGA_VSYNC_NEG,
	RESULT
);


//=======================================================
//  PORT declarations
//=======================================================
input	[7:0]	PIXEL_IN;
input			CLK;
input [9:0]	VGA_PIXEL_X;
input	[9:0]	VGA_PIXEL_Y;
input			VGA_VSYNC_NEG;

output reg [2:0] RESULT;

reg [15:0] BLUECOUNTTOP = 0;
reg [15:0] REDCOUNTTOP = 0;
reg [15:0] BLUECOUNTMID = 0;
reg [15:0] REDCOUNTMID = 0;
reg [15:0] BLUECOUNTBOTTOM = 0;
reg [15:0] REDCOUNTBOTTOM = 0;
reg [15:0] REDCOUNTTEMPTOP = 0;
reg [15:0] BLUECOUNTTEMPTOP = 0;
reg [15:0] REDCOUNTTEMPMID = 0;
reg [15:0] BLUECOUNTTEMPMID = 0;
reg [15:0] REDCOUNTTEMPBOTTOM = 0;
reg [15:0] BLUECOUNTTEMPBOTTOM = 0;

always @ (posedge CLK, negedge VGA_VSYNC_NEG) begin
		if (!VGA_VSYNC_NEG) begin
			if ((BLUECOUNTTEMPTOP+BLUECOUNTTEMPBOTTOM+BLUECOUNTTEMPMID) > (REDCOUNTTEMPTOP+REDCOUNTBOTTOM+REDCOUNTTEMPMID) && (BLUECOUNTTEMPTOP+BLUECOUNTTEMPBOTTOM+BLUECOUNTTEMPMID) > 16'd10000) begin //17000 is arbitrary, can change
				if (BLUECOUNTTEMPTOP<BLUECOUNTTEMPMID && BLUECOUNTTEMPMID<BLUECOUNTTEMPBOTTOM) begin //&& BLUECOUNTTEMPTOP<BLUECOUNTTEMPBOTTOM 
					RESULT = 3'b001; //blue triangle
				end
				else if (BLUECOUNTTEMPTOP<BLUECOUNTTEMPMID && BLUECOUNTTEMPMID>BLUECOUNTTEMPBOTTOM && (BLUECOUNTTEMPBOTTOM<=(BLUECOUNTTEMPTOP+20) && BLUECOUNTTEMPBOTTOM>=(BLUECOUNTTEMPTOP-20))) begin
					RESULT = 3'b010; //blue diamond
				end
				else begin
					RESULT = 3'b011; //blue square
				end
			end
			else if ((REDCOUNTTEMPTOP+REDCOUNTTEMPBOTTOM+REDCOUNTTEMPMID) > (BLUECOUNTTEMPTOP+BLUECOUNTBOTTOM+BLUECOUNTTEMPMID) && (REDCOUNTTEMPTOP+REDCOUNTTEMPBOTTOM+REDCOUNTTEMPMID) > 16'd10000) begin //17000 is arbitrary, can change
				if (REDCOUNTTEMPTOP<REDCOUNTTEMPMID && REDCOUNTTEMPMID>REDCOUNTTEMPBOTTOM) begin //&& REDCOUNTTEMPTOP<REDCOUNTTEMPBOTTOM 
					RESULT = 3'b100; //red triangle
				end
				else if (REDCOUNTTEMPTOP<REDCOUNTTEMPMID && REDCOUNTTEMPMID>REDCOUNTTEMPBOTTOM && (REDCOUNTTEMPBOTTOM<=(REDCOUNTTEMPTOP+20) && REDCOUNTTEMPBOTTOM>=(REDCOUNTTEMPTOP-20))) begin
					RESULT = 3'b101; //red diamond
				end
				else begin
					RESULT = 3'b110; //red square
				end
			end
			else begin
				RESULT = 3'b000; //no color detected
			end
			BLUECOUNTTOP = 0;
			REDCOUNTTOP = 0;
			BLUECOUNTMID = 0;
			REDCOUNTMID = 0;
			BLUECOUNTBOTTOM = 0;
			REDCOUNTBOTTOM = 0;
		end
		else begin
			RESULT = RESULT;
			if (VGA_PIXEL_Y >= 10'd30 && VGA_PIXEL_Y <= 10'd59) begin
				if (PIXEL_IN[7:6] > PIXEL_IN[1:0] && PIXEL_IN[7:6] > PIXEL_IN[4:3]) begin
					REDCOUNTTOP = REDCOUNTTOP + 1'b1;
				end
				else if (PIXEL_IN[1:0] > PIXEL_IN[7:6] && PIXEL_IN[1:0] > PIXEL_IN[4:3]) begin
					BLUECOUNTTOP = BLUECOUNTTOP + 1'b1;
				end
				REDCOUNTTEMPTOP = REDCOUNTTOP;
				BLUECOUNTTEMPTOP = BLUECOUNTTOP;
			end
			else if (VGA_PIXEL_Y >= 10'd60 && VGA_PIXEL_Y <= 10'd89) begin
				if (PIXEL_IN[7:6] > PIXEL_IN[1:0] && PIXEL_IN[7:6] > PIXEL_IN[4:3]) begin
					REDCOUNTMID = REDCOUNTMID + 1'b1;
				end
				else if (PIXEL_IN[1:0] > PIXEL_IN[7:6] && PIXEL_IN[1:0] > PIXEL_IN[4:3]) begin
					BLUECOUNTMID = BLUECOUNTMID + 1'b1;
				end
				REDCOUNTTEMPMID = REDCOUNTMID;
				BLUECOUNTTEMPMID = BLUECOUNTMID;
			end
			else if (VGA_PIXEL_Y >= 10'd90 && VGA_PIXEL_Y <= 10'd119) begin
				if (PIXEL_IN[7:6] > PIXEL_IN[1:0] && PIXEL_IN[7:6] > PIXEL_IN[4:3]) begin
					REDCOUNTBOTTOM = REDCOUNTBOTTOM + 1'b1;
				end
				else if (PIXEL_IN[1:0] > PIXEL_IN[7:6] && PIXEL_IN[1:0] > PIXEL_IN[4:3]) begin
					BLUECOUNTBOTTOM = BLUECOUNTBOTTOM + 1'b1;
				end
				REDCOUNTTEMPBOTTOM = REDCOUNTBOTTOM;
				BLUECOUNTTEMPBOTTOM = BLUECOUNTBOTTOM;
			end
		end
end


endmodule